
reg dev_state; // 0- это init 1- это работа по установке угла
reg [7:0] angle_target; //целевой
reg [7:0] angle_current; //текущий

endmodule
