module RELAY1 (input A, input B, output Q);
assign Q = A & B; 
endmodule